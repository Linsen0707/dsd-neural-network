--beginning case
s(0)=a(0)AND b(0)

--end case
s(15)=a(7)AND b(7)

--normal case
int p=cnt-1;
for(int q=0; q<cnt; q++) {
	--generate adders
	Adder: FullAdder
		port map(a(p),b(
	--decrement counter
	p=p-1;
}